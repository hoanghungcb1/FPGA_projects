library verilog;
use verilog.vl_types.all;
entity wrapper_9_vlg_check_tst is
    port(
        P               : in     vl_logic_vector(15 downto 0);
        sampler_rx      : in     vl_logic
    );
end wrapper_9_vlg_check_tst;
