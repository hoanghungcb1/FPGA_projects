library verilog;
use verilog.vl_types.all;
entity wrapper_9_vlg_vec_tst is
end wrapper_9_vlg_vec_tst;
