library verilog;
use verilog.vl_types.all;
entity wrapper_8_vlg_vec_tst is
end wrapper_8_vlg_vec_tst;
